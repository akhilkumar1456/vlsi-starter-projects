module hello;
  initial begin
    $display("--- Hello World! Compilation Test Successful ---");
    $finish;
  end
endmodule