// MUX2x1.v
module MUX2x1 (
    input D0,   // Check spelling: D0, D1, S
    input D1,   
    input S,    
    output Y    // Check spelling: Y
);
// ... logic here ...
endmodule